module top_module (
    input clk,
    input enable,
    input S,
    input A, B, C,
    output Z ); 

reg [7:0] Q;
always @(posedge clk ) begin
    if (enable) begin
        Q <= {Q[7:1],S};
    end else begin
        Q <= Q;
    end
end

assign Z = Q[{A,B,C}]; 
endmodule